`define DATA_WIDTH 4

`define MODE0   4'd0    // add
`define MODE1   4'd1    // subtract
`define MODE2   4'd2    // multiply
`define MODE3   4'd3    // divide
`define MODE4   4'd4    // left shift logical
`define MODE5   4'd5    // right shift logical
`define MODE6   4'd6    // rotate left
`define MODE7   4'd7    // rotate right
`define MODE8   4'd8    // logical and
`define MODE9   4'd9    // logical or
`define MODE10  4'd10   // logical xor
`define MODE11  4'd11   // logical nand
`define MODE12  4'd12   // logical nor
`define MODE13  4'd13   // logical xnor
`define MODE14  4'd14   // greater comparison
`define MODE15  4'd15   // equal comparison
